// COMMIT: modbus串口服务模块
// DSC:
// 	接收总线上的数据，发出数据和数据有效标志

module mbUartR(
    port_list
);
    
endmodule
// COMMIT: modbus串口服务模块
// DSC:
// 	接收数据和数据有效标志，通过串口发出，返回发送完成标志

module mbUartT(
    port_list
);
    
endmodule
// COMMIT: 传感器接收数据汇总模块
// DSC:
// 	接收来自各个串口接收模块的消息
// 	发送给数据缓存模块

module rxcomb(
	input			sys_clk,
	input			sys_rst,	
	
	
	
);



endmodule
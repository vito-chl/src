// COMMIT: 传感器发送数据汇总模块
// DSC:
// 	接收配置命令，控制一段时间内发送传感器数据请求命令
// 	发送给各种形式的发送模块

module txcomb(
	input			sys_clk,
	input			sys_rst,
	
	
);




endmodule
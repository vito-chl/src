module tranbus(
	
);




endmodule
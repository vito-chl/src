// COMMIT: 总线数据接收解析模块
// DSC:
// 	解析来自总线的数据，进行相应处理，并发送给总线数据生成模块
//	或者发送给传感器命令模块

module rxana(
	input			sys_clk,
	input			sys_rst,
	
	// 消息接收模块接收到的消息
	input			rx_flag,// 接收数据完成的标志
	input	[7:0]	rx_data,// 接收的数据
	
	// 总线数据生成模块
	output 	[x:0]	ret_cmd, // 返回命令
	output			ret_cmd_flg, // 返回命令有效标志
	
	// 传感器命令模块
	output	[x:0]	sen_cmd, // 发送的命令
	output	[x:0]	data	// 发送的数据
);

//*****************************  接口协议  *****************************
// * 数据<rx_data>准备好，同时给接收标志<rx_flag>一个周期的高电平
// * 命令<ret_cmd>会提前准备好，同时有效标志<ret_cmd_flg> 
//   会给一个周期的高电平
// * 数据<data>会提前准备好，同时发送一个周期命令<sen_cmd>
//**********************************************************************

//*****************************  mianStaM  *****************************
// * 
//**********************************************************************
reg []


endmodule